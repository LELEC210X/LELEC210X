// (C) 2001-2018 Intel Corporation. All rights reserved.
<<<<<<< refs/remotes/upstream/main
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
=======
// Your use of Intel Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions, and any output
// files from any of the foregoing (including device programming or simulation
// files), and any associated documentation or information are expressly subject
// to the terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other applicable
// license agreement, including, without limitation, that your use is for the
// sole purpose of programming logic devices manufactured by Intel and sold by
// Intel or its authorized distributors.  Please refer to the applicable
>>>>>>> Revert "enlever le chain de argu"
// agreement for further details.



<<<<<<< refs/remotes/upstream/main
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
=======
// Your use of Altera Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions, and any output
// files any of the foregoing (including device programming or simulation
// files), and any associated documentation or information are expressly subject
// to the terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other applicable
// license agreement, including, without limitation, that your use is for the
// sole purpose of programming logic devices manufactured by Altera and sold by
// Altera or its authorized distributors.  Please refer to the applicable
>>>>>>> Revert "enlever le chain de argu"
// agreement for further details.


// $Id: //acds/rel/18.1std/ip/merlin/altera_merlin_router/altera_merlin_router.sv.terp#1 $
// $Revision: #1 $
// $Date: 2018/07/18 $
// $Author: psgswbuild $

// -------------------------------------------------------
// Merlin Router
//
<<<<<<< refs/remotes/upstream/main
// Asserts the appropriate one-hot encoded channel based on 
=======
// Asserts the appropriate one-hot encoded channel based on
>>>>>>> Revert "enlever le chain de argu"
// either (a) the address or (b) the dest id. The DECODER_TYPE
// parameter controls this behaviour. 0 means address decoder,
// 1 means dest id decoder.
//
// In the case of (a), it also sets the destination id.
// -------------------------------------------------------

`timescale 1 ns / 1 ns

module lms_ctr_mm_interconnect_0_router_default_decode
  #(
     parameter DEFAULT_CHANNEL = 5,
               DEFAULT_WR_CHANNEL = -1,
               DEFAULT_RD_CHANNEL = -1,
<<<<<<< refs/remotes/upstream/main
               DEFAULT_DESTID = 10 
=======
               DEFAULT_DESTID = 10
>>>>>>> Revert "enlever le chain de argu"
   )
  (output [89 - 86 : 0] default_destination_id,
   output [15-1 : 0] default_wr_channel,
   output [15-1 : 0] default_rd_channel,
   output [15-1 : 0] default_src_channel
  );

<<<<<<< refs/remotes/upstream/main
  assign default_destination_id = 
=======
  assign default_destination_id =
>>>>>>> Revert "enlever le chain de argu"
    DEFAULT_DESTID[89 - 86 : 0];

  generate
    if (DEFAULT_CHANNEL == -1) begin : no_default_channel_assignment
      assign default_src_channel = '0;
    end
    else begin : default_channel_assignment
      assign default_src_channel = 15'b1 << DEFAULT_CHANNEL;
    end
  endgenerate

  generate
    if (DEFAULT_RD_CHANNEL == -1) begin : no_default_rw_channel_assignment
      assign default_wr_channel = '0;
      assign default_rd_channel = '0;
    end
    else begin : default_rw_channel_assignment
      assign default_wr_channel = 15'b1 << DEFAULT_WR_CHANNEL;
      assign default_rd_channel = 15'b1 << DEFAULT_RD_CHANNEL;
    end
  endgenerate

endmodule


module lms_ctr_mm_interconnect_0_router
(
    // -------------------
    // Clock & Reset
    // -------------------
    input clk,
    input reset,

    // -------------------
    // Command Sink (Input)
    // -------------------
    input                       sink_valid,
    input  [103-1 : 0]    sink_data,
    input                       sink_startofpacket,
    input                       sink_endofpacket,
    output                      sink_ready,

    // -------------------
    // Command Source (Output)
    // -------------------
    output                          src_valid,
    output reg [103-1    : 0] src_data,
    output reg [15-1 : 0] src_channel,
    output                          src_startofpacket,
    output                          src_endofpacket,
    input                           src_ready
);

    // -------------------------------------------------------
    // Local parameters and variables
    // -------------------------------------------------------
    localparam PKT_ADDR_H = 57;
    localparam PKT_ADDR_L = 36;
    localparam PKT_DEST_ID_H = 89;
    localparam PKT_DEST_ID_L = 86;
    localparam PKT_PROTECTION_H = 93;
    localparam PKT_PROTECTION_L = 91;
    localparam ST_DATA_W = 103;
    localparam ST_CHANNEL_W = 15;
    localparam DECODER_TYPE = 0;

    localparam PKT_TRANS_WRITE = 60;
    localparam PKT_TRANS_READ  = 61;

    localparam PKT_ADDR_W = PKT_ADDR_H-PKT_ADDR_L + 1;
    localparam PKT_DEST_ID_W = PKT_DEST_ID_H-PKT_DEST_ID_L + 1;



    // -------------------------------------------------------
    // Figure out the number of bits to mask off for each slave span
    // during address decoding
    // -------------------------------------------------------
<<<<<<< refs/remotes/upstream/main
    localparam PAD0 = log2ceil(64'h200000 - 64'h100000); 
    localparam PAD1 = log2ceil(64'h201000 - 64'h200000); 
    localparam PAD2 = log2ceil(64'h202000 - 64'h201800); 
    localparam PAD3 = log2ceil(64'h202020 - 64'h202000); 
    localparam PAD4 = log2ceil(64'h202040 - 64'h202020); 
    localparam PAD5 = log2ceil(64'h202060 - 64'h202040); 
    localparam PAD6 = log2ceil(64'h202080 - 64'h202060); 
    localparam PAD7 = log2ceil(64'h2020a0 - 64'h202080); 
    localparam PAD8 = log2ceil(64'h2020c0 - 64'h2020a0); 
    localparam PAD9 = log2ceil(64'h2020e0 - 64'h2020c0); 
    localparam PAD10 = log2ceil(64'h2020f0 - 64'h2020e0); 
    localparam PAD11 = log2ceil(64'h202100 - 64'h2020f0); 
    localparam PAD12 = log2ceil(64'h202110 - 64'h202100); 
    localparam PAD13 = log2ceil(64'h202118 - 64'h202110); 
    localparam PAD14 = log2ceil(64'h202120 - 64'h202118); 
=======
    localparam PAD0 = log2ceil(64'h200000 - 64'h100000);
    localparam PAD1 = log2ceil(64'h201000 - 64'h200000);
    localparam PAD2 = log2ceil(64'h202000 - 64'h201800);
    localparam PAD3 = log2ceil(64'h202020 - 64'h202000);
    localparam PAD4 = log2ceil(64'h202040 - 64'h202020);
    localparam PAD5 = log2ceil(64'h202060 - 64'h202040);
    localparam PAD6 = log2ceil(64'h202080 - 64'h202060);
    localparam PAD7 = log2ceil(64'h2020a0 - 64'h202080);
    localparam PAD8 = log2ceil(64'h2020c0 - 64'h2020a0);
    localparam PAD9 = log2ceil(64'h2020e0 - 64'h2020c0);
    localparam PAD10 = log2ceil(64'h2020f0 - 64'h2020e0);
    localparam PAD11 = log2ceil(64'h202100 - 64'h2020f0);
    localparam PAD12 = log2ceil(64'h202110 - 64'h202100);
    localparam PAD13 = log2ceil(64'h202118 - 64'h202110);
    localparam PAD14 = log2ceil(64'h202120 - 64'h202118);
>>>>>>> Revert "enlever le chain de argu"
    // -------------------------------------------------------
    // Work out which address bits are significant based on the
    // address range of the slaves. If the required width is too
    // large or too small, we use the address field width instead.
    // -------------------------------------------------------
    localparam ADDR_RANGE = 64'h202120;
    localparam RANGE_ADDR_WIDTH = log2ceil(ADDR_RANGE);
    localparam OPTIMIZED_ADDR_H = (RANGE_ADDR_WIDTH > PKT_ADDR_W) ||
                                  (RANGE_ADDR_WIDTH == 0) ?
                                        PKT_ADDR_H :
                                        PKT_ADDR_L + RANGE_ADDR_WIDTH - 1;

    localparam RG = RANGE_ADDR_WIDTH-1;
    localparam REAL_ADDRESS_RANGE = OPTIMIZED_ADDR_H - PKT_ADDR_L;

      reg [PKT_ADDR_W-1 : 0] address;
      always @* begin
        address = {PKT_ADDR_W{1'b0}};
        address [REAL_ADDRESS_RANGE:0] = sink_data[OPTIMIZED_ADDR_H : PKT_ADDR_L];
<<<<<<< refs/remotes/upstream/main
      end   
=======
      end
>>>>>>> Revert "enlever le chain de argu"

    // -------------------------------------------------------
    // Pass almost everything through, untouched
    // -------------------------------------------------------
    assign sink_ready        = src_ready;
    assign src_valid         = sink_valid;
    assign src_startofpacket = sink_startofpacket;
    assign src_endofpacket   = sink_endofpacket;
    wire [PKT_DEST_ID_W-1:0] default_destid;
    wire [15-1 : 0] default_src_channel;




    // -------------------------------------------------------
    // Write and read transaction signals
    // -------------------------------------------------------
    wire read_transaction;
    assign read_transaction  = sink_data[PKT_TRANS_READ];


    lms_ctr_mm_interconnect_0_router_default_decode the_default_decode(
      .default_destination_id (default_destid),
      .default_wr_channel   (),
      .default_rd_channel   (),
      .default_src_channel  (default_src_channel)
    );

    always @* begin
        src_data    = sink_data;
        src_channel = default_src_channel;
        src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = default_destid;

        // --------------------------------------------------
        // Address Decoder
        // Sets the channel and destination ID based on the address
        // --------------------------------------------------

    // ( 0x100000 .. 0x200000 )
    if ( {address[RG:PAD0],{PAD0{1'b0}}} == 22'h100000   ) begin
            src_channel = 15'b000000000100000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 10;
    end

    // ( 0x200000 .. 0x201000 )
    if ( {address[RG:PAD1],{PAD1{1'b0}}} == 22'h200000   ) begin
            src_channel = 15'b000100000000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 11;
    end

    // ( 0x201800 .. 0x202000 )
    if ( {address[RG:PAD2],{PAD2{1'b0}}} == 22'h201800   ) begin
            src_channel = 15'b000000001000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 8;
    end

    // ( 0x202000 .. 0x202020 )
    if ( {address[RG:PAD3],{PAD3{1'b0}}} == 22'h202000   ) begin
            src_channel = 15'b100000000000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 3;
    end

    // ( 0x202020 .. 0x202040 )
    if ( {address[RG:PAD4],{PAD4{1'b0}}} == 22'h202020   ) begin
            src_channel = 15'b010000000000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 1;
    end

    // ( 0x202040 .. 0x202060 )
    if ( {address[RG:PAD5],{PAD5{1'b0}}} == 22'h202040   ) begin
            src_channel = 15'b001000000000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 4;
    end

    // ( 0x202060 .. 0x202080 )
    if ( {address[RG:PAD6],{PAD6{1'b0}}} == 22'h202060   ) begin
            src_channel = 15'b000010000000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 7;
    end

    // ( 0x202080 .. 0x2020a0 )
    if ( {address[RG:PAD7],{PAD7{1'b0}}} == 22'h202080   ) begin
            src_channel = 15'b000001000000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 14;
    end

    // ( 0x2020a0 .. 0x2020c0 )
    if ( {address[RG:PAD8],{PAD8{1'b0}}} == 22'h2020a0   ) begin
            src_channel = 15'b000000000000100;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 5;
    end

    // ( 0x2020c0 .. 0x2020e0 )
    if ( {address[RG:PAD9],{PAD9{1'b0}}} == 22'h2020c0   ) begin
            src_channel = 15'b000000000000001;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 2;
    end

    // ( 0x2020e0 .. 0x2020f0 )
    if ( {address[RG:PAD10],{PAD10{1'b0}}} == 22'h2020e0   ) begin
            src_channel = 15'b000000100000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 6;
    end

    // ( 0x2020f0 .. 0x202100 )
    if ( {address[RG:PAD11],{PAD11{1'b0}}} == 22'h2020f0  && read_transaction  ) begin
            src_channel = 15'b000000010000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 12;
    end

    // ( 0x202100 .. 0x202110 )
    if ( {address[RG:PAD12],{PAD12{1'b0}}} == 22'h202100   ) begin
            src_channel = 15'b000000000000010;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 0;
    end

    // ( 0x202110 .. 0x202118 )
    if ( {address[RG:PAD13],{PAD13{1'b0}}} == 22'h202110   ) begin
            src_channel = 15'b000000000010000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 9;
    end

    // ( 0x202118 .. 0x202120 )
    if ( {address[RG:PAD14],{PAD14{1'b0}}} == 22'h202118  && read_transaction  ) begin
            src_channel = 15'b000000000001000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 13;
    end

end


    // --------------------------------------------------
    // Ceil(log2()) function
    // --------------------------------------------------
    function integer log2ceil;
        input reg[65:0] val;
        reg [65:0] i;

        begin
            i = 1;
            log2ceil = 0;

            while (i < val) begin
                log2ceil = log2ceil + 1;
                i = i << 1;
            end
        end
    endfunction

endmodule
<<<<<<< refs/remotes/upstream/main


=======
>>>>>>> Revert "enlever le chain de argu"
