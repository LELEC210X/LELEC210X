// lms_ctr.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module lms_ctr (
		input  wire        clk_clk,                                 //                              clk.clk
		input  wire        dac_spi_ext_MISO,                        //                      dac_spi_ext.MISO
		output wire        dac_spi_ext_MOSI,                        //                                 .MOSI
		output wire        dac_spi_ext_SCLK,                        //                                 .SCLK
		output wire        dac_spi_ext_SS_n,                        //                                 .SS_n
		input  wire [31:0] exfifo_if_d_export,                      //                      exfifo_if_d.export
		output wire        exfifo_if_rd_export,                     //                     exfifo_if_rd.export
		input  wire        exfifo_if_rdempty_export,                //                exfifo_if_rdempty.export
		output wire [31:0] exfifo_of_d_export,                      //                      exfifo_of_d.export
		output wire        exfifo_of_wr_export,                     //                     exfifo_of_wr.export
		input  wire        exfifo_of_wrfull_export,                 //                 exfifo_of_wrfull.export
		output wire        exfifo_rst_export,                       //                       exfifo_rst.export
		input  wire        flash_spi_MISO,                          //                        flash_spi.MISO
		output wire        flash_spi_MOSI,                          //                                 .MOSI
		output wire        flash_spi_SCLK,                          //                                 .SCLK
		output wire        flash_spi_SS_n,                          //                                 .SS_n
		input  wire        fpga_spi_ext_MISO,                       //                     fpga_spi_ext.MISO
		output wire        fpga_spi_ext_MOSI,                       //                                 .MOSI
		output wire        fpga_spi_ext_SCLK,                       //                                 .SCLK
		output wire [1:0]  fpga_spi_ext_SS_n,                       //                                 .SS_n
		inout  wire        i2c_scl_export,                          //                          i2c_scl.export
		inout  wire        i2c_sda_export,                          //                          i2c_sda.export
		output wire [7:0]  leds_external_connection_export,         //         leds_external_connection.export
		output wire [3:0]  lms_ctr_gpio_external_connection_export, // lms_ctr_gpio_external_connection.export
		input  wire [7:0]  switch_external_connection_export,       //       switch_external_connection.export
		input  wire        uart_external_connection_rxd,            //         uart_external_connection.rxd
		output wire        uart_external_connection_txd             //                                 .txd
	);

	wire         nios2_cpu_debug_reset_request_reset;                                         // nios2_cpu:debug_reset_request -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire         nios2_cpu_custom_instruction_master_readra;                                  // nios2_cpu:D_ci_readra -> nios2_cpu_custom_instruction_master_translator:ci_slave_readra
	wire   [4:0] nios2_cpu_custom_instruction_master_a;                                       // nios2_cpu:D_ci_a -> nios2_cpu_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] nios2_cpu_custom_instruction_master_b;                                       // nios2_cpu:D_ci_b -> nios2_cpu_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios2_cpu_custom_instruction_master_c;                                       // nios2_cpu:D_ci_c -> nios2_cpu_custom_instruction_master_translator:ci_slave_c
	wire         nios2_cpu_custom_instruction_master_readrb;                                  // nios2_cpu:D_ci_readrb -> nios2_cpu_custom_instruction_master_translator:ci_slave_readrb
	wire  [31:0] nios2_cpu_custom_instruction_master_ipending;                                // nios2_cpu:W_ci_ipending -> nios2_cpu_custom_instruction_master_translator:ci_slave_ipending
	wire   [7:0] nios2_cpu_custom_instruction_master_n;                                       // nios2_cpu:D_ci_n -> nios2_cpu_custom_instruction_master_translator:ci_slave_n
	wire  [31:0] nios2_cpu_custom_instruction_master_result;                                  // nios2_cpu_custom_instruction_master_translator:ci_slave_result -> nios2_cpu:E_ci_result
	wire         nios2_cpu_custom_instruction_master_estatus;                                 // nios2_cpu:W_ci_estatus -> nios2_cpu_custom_instruction_master_translator:ci_slave_estatus
	wire  [31:0] nios2_cpu_custom_instruction_master_datab;                                   // nios2_cpu:E_ci_datab -> nios2_cpu_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] nios2_cpu_custom_instruction_master_dataa;                                   // nios2_cpu:E_ci_dataa -> nios2_cpu_custom_instruction_master_translator:ci_slave_dataa
	wire         nios2_cpu_custom_instruction_master_writerc;                                 // nios2_cpu:D_ci_writerc -> nios2_cpu_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_result;        // nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_result -> nios2_cpu_custom_instruction_master_translator:comb_ci_master_result
	wire         nios2_cpu_custom_instruction_master_translator_comb_ci_master_readra;        // nios2_cpu_custom_instruction_master_translator:comb_ci_master_readra -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_a;             // nios2_cpu_custom_instruction_master_translator:comb_ci_master_a -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_b;             // nios2_cpu_custom_instruction_master_translator:comb_ci_master_b -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         nios2_cpu_custom_instruction_master_translator_comb_ci_master_readrb;        // nios2_cpu_custom_instruction_master_translator:comb_ci_master_readrb -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_c;             // nios2_cpu_custom_instruction_master_translator:comb_ci_master_c -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         nios2_cpu_custom_instruction_master_translator_comb_ci_master_estatus;       // nios2_cpu_custom_instruction_master_translator:comb_ci_master_estatus -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_ipending;      // nios2_cpu_custom_instruction_master_translator:comb_ci_master_ipending -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_datab;         // nios2_cpu_custom_instruction_master_translator:comb_ci_master_datab -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_dataa;         // nios2_cpu_custom_instruction_master_translator:comb_ci_master_dataa -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         nios2_cpu_custom_instruction_master_translator_comb_ci_master_writerc;       // nios2_cpu_custom_instruction_master_translator:comb_ci_master_writerc -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_n;             // nios2_cpu_custom_instruction_master_translator:comb_ci_master_n -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_result;         // nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_result -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readra;         // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_readra -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_a;              // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_a -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_b;              // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_b -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb;         // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_readrb -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_c;              // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_c -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus;        // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_estatus -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending;       // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_ipending -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_datab;          // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_datab -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa;          // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_dataa -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc;        // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_writerc -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_n;              // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_n -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_result; // nios_custom_instr_bitswap_0:result -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab;  // nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_master_datab -> nios_custom_instr_bitswap_0:datab
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa;  // nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> nios_custom_instr_bitswap_0:dataa
	wire  [31:0] nios2_cpu_data_master_readdata;                                              // mm_interconnect_0:nios2_cpu_data_master_readdata -> nios2_cpu:d_readdata
	wire         nios2_cpu_data_master_waitrequest;                                           // mm_interconnect_0:nios2_cpu_data_master_waitrequest -> nios2_cpu:d_waitrequest
	wire         nios2_cpu_data_master_debugaccess;                                           // nios2_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_cpu_data_master_debugaccess
	wire  [21:0] nios2_cpu_data_master_address;                                               // nios2_cpu:d_address -> mm_interconnect_0:nios2_cpu_data_master_address
	wire   [3:0] nios2_cpu_data_master_byteenable;                                            // nios2_cpu:d_byteenable -> mm_interconnect_0:nios2_cpu_data_master_byteenable
	wire         nios2_cpu_data_master_read;                                                  // nios2_cpu:d_read -> mm_interconnect_0:nios2_cpu_data_master_read
	wire         nios2_cpu_data_master_write;                                                 // nios2_cpu:d_write -> mm_interconnect_0:nios2_cpu_data_master_write
	wire  [31:0] nios2_cpu_data_master_writedata;                                             // nios2_cpu:d_writedata -> mm_interconnect_0:nios2_cpu_data_master_writedata
	wire  [31:0] nios2_cpu_instruction_master_readdata;                                       // mm_interconnect_0:nios2_cpu_instruction_master_readdata -> nios2_cpu:i_readdata
	wire         nios2_cpu_instruction_master_waitrequest;                                    // mm_interconnect_0:nios2_cpu_instruction_master_waitrequest -> nios2_cpu:i_waitrequest
	wire  [21:0] nios2_cpu_instruction_master_address;                                        // nios2_cpu:i_address -> mm_interconnect_0:nios2_cpu_instruction_master_address
	wire         nios2_cpu_instruction_master_read;                                           // nios2_cpu:i_read -> mm_interconnect_0:nios2_cpu_instruction_master_read
	wire  [31:0] mm_interconnect_0_dual_boot_0_avalon_readdata;                               // dual_boot_0:avmm_rcv_readdata -> mm_interconnect_0:dual_boot_0_avalon_readdata
	wire   [2:0] mm_interconnect_0_dual_boot_0_avalon_address;                                // mm_interconnect_0:dual_boot_0_avalon_address -> dual_boot_0:avmm_rcv_address
	wire         mm_interconnect_0_dual_boot_0_avalon_read;                                   // mm_interconnect_0:dual_boot_0_avalon_read -> dual_boot_0:avmm_rcv_read
	wire         mm_interconnect_0_dual_boot_0_avalon_write;                                  // mm_interconnect_0:dual_boot_0_avalon_write -> dual_boot_0:avmm_rcv_write
	wire  [31:0] mm_interconnect_0_dual_boot_0_avalon_writedata;                              // mm_interconnect_0:dual_boot_0_avalon_writedata -> dual_boot_0:avmm_rcv_writedata
	wire         mm_interconnect_0_av_fifo_int_0_avalon_slave_0_chipselect;                   // mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_chipselect -> Av_FIFO_Int_0:chipselect
	wire  [31:0] mm_interconnect_0_av_fifo_int_0_avalon_slave_0_readdata;                     // Av_FIFO_Int_0:readdata -> mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_av_fifo_int_0_avalon_slave_0_address;                      // mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_address -> Av_FIFO_Int_0:address
	wire         mm_interconnect_0_av_fifo_int_0_avalon_slave_0_read;                         // mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_read -> Av_FIFO_Int_0:read
	wire         mm_interconnect_0_av_fifo_int_0_avalon_slave_0_write;                        // mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_write -> Av_FIFO_Int_0:write
	wire  [31:0] mm_interconnect_0_av_fifo_int_0_avalon_slave_0_writedata;                    // mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_writedata -> Av_FIFO_Int_0:writedata
	wire         mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect;                 // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_chipselect -> i2c_opencores_0:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata;                   // i2c_opencores_0:wb_dat_o -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_i2c_opencores_0_avalon_slave_0_waitrequest;                // i2c_opencores_0:wb_ack_o -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address;                    // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_address -> i2c_opencores_0:wb_adr_i
	wire         mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write;                      // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_write -> i2c_opencores_0:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata;                  // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_writedata -> i2c_opencores_0:wb_dat_i
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;                       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;                        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_readdata;                               // onchip_flash_0:avmm_csr_readdata -> mm_interconnect_0:onchip_flash_0_csr_readdata
	wire   [0:0] mm_interconnect_0_onchip_flash_0_csr_address;                                // mm_interconnect_0:onchip_flash_0_csr_address -> onchip_flash_0:avmm_csr_addr
	wire         mm_interconnect_0_onchip_flash_0_csr_read;                                   // mm_interconnect_0:onchip_flash_0_csr_read -> onchip_flash_0:avmm_csr_read
	wire         mm_interconnect_0_onchip_flash_0_csr_write;                                  // mm_interconnect_0:onchip_flash_0_csr_write -> onchip_flash_0:avmm_csr_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_writedata;                              // mm_interconnect_0:onchip_flash_0_csr_writedata -> onchip_flash_0:avmm_csr_writedata
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_readdata;                              // onchip_flash_0:avmm_data_readdata -> mm_interconnect_0:onchip_flash_0_data_readdata
	wire         mm_interconnect_0_onchip_flash_0_data_waitrequest;                           // onchip_flash_0:avmm_data_waitrequest -> mm_interconnect_0:onchip_flash_0_data_waitrequest
	wire  [17:0] mm_interconnect_0_onchip_flash_0_data_address;                               // mm_interconnect_0:onchip_flash_0_data_address -> onchip_flash_0:avmm_data_addr
	wire         mm_interconnect_0_onchip_flash_0_data_read;                                  // mm_interconnect_0:onchip_flash_0_data_read -> onchip_flash_0:avmm_data_read
	wire         mm_interconnect_0_onchip_flash_0_data_readdatavalid;                         // onchip_flash_0:avmm_data_readdatavalid -> mm_interconnect_0:onchip_flash_0_data_readdatavalid
	wire         mm_interconnect_0_onchip_flash_0_data_write;                                 // mm_interconnect_0:onchip_flash_0_data_write -> onchip_flash_0:avmm_data_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_writedata;                             // mm_interconnect_0:onchip_flash_0_data_writedata -> onchip_flash_0:avmm_data_writedata
	wire   [3:0] mm_interconnect_0_onchip_flash_0_data_burstcount;                            // mm_interconnect_0:onchip_flash_0_data_burstcount -> onchip_flash_0:avmm_data_burstcount
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata;                        // nios2_cpu:debug_mem_slave_readdata -> mm_interconnect_0:nios2_cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest;                     // nios2_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess;                     // mm_interconnect_0:nios2_cpu_debug_mem_slave_debugaccess -> nios2_cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_address;                         // mm_interconnect_0:nios2_cpu_debug_mem_slave_address -> nios2_cpu:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_read;                            // mm_interconnect_0:nios2_cpu_debug_mem_slave_read -> nios2_cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable;                      // mm_interconnect_0:nios2_cpu_debug_mem_slave_byteenable -> nios2_cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_write;                           // mm_interconnect_0:nios2_cpu_debug_mem_slave_write -> nios2_cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata;                       // mm_interconnect_0:nios2_cpu_debug_mem_slave_writedata -> nios2_cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_switch_s1_readdata;                                        // switch:readdata -> mm_interconnect_0:switch_s1_readdata
	wire   [1:0] mm_interconnect_0_switch_s1_address;                                         // mm_interconnect_0:switch_s1_address -> switch:address
	wire         mm_interconnect_0_leds_s1_chipselect;                                        // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                          // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                           // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_write;                                             // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                         // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire         mm_interconnect_0_uart_s1_chipselect;                                        // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                                          // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                                           // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_read;                                              // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;                                     // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                                             // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                                         // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire         mm_interconnect_0_lms_ctr_gpio_s1_chipselect;                                // mm_interconnect_0:lms_ctr_gpio_s1_chipselect -> lms_ctr_gpio:chipselect
	wire  [31:0] mm_interconnect_0_lms_ctr_gpio_s1_readdata;                                  // lms_ctr_gpio:readdata -> mm_interconnect_0:lms_ctr_gpio_s1_readdata
	wire   [2:0] mm_interconnect_0_lms_ctr_gpio_s1_address;                                   // mm_interconnect_0:lms_ctr_gpio_s1_address -> lms_ctr_gpio:address
	wire         mm_interconnect_0_lms_ctr_gpio_s1_write;                                     // mm_interconnect_0:lms_ctr_gpio_s1_write -> lms_ctr_gpio:write_n
	wire  [31:0] mm_interconnect_0_lms_ctr_gpio_s1_writedata;                                 // mm_interconnect_0:lms_ctr_gpio_s1_writedata -> lms_ctr_gpio:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;                               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_fpga_spi_spi_control_port_chipselect;                      // mm_interconnect_0:fpga_spi_spi_control_port_chipselect -> fpga_spi:spi_select
	wire  [15:0] mm_interconnect_0_fpga_spi_spi_control_port_readdata;                        // fpga_spi:data_to_cpu -> mm_interconnect_0:fpga_spi_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_fpga_spi_spi_control_port_address;                         // mm_interconnect_0:fpga_spi_spi_control_port_address -> fpga_spi:mem_addr
	wire         mm_interconnect_0_fpga_spi_spi_control_port_read;                            // mm_interconnect_0:fpga_spi_spi_control_port_read -> fpga_spi:read_n
	wire         mm_interconnect_0_fpga_spi_spi_control_port_write;                           // mm_interconnect_0:fpga_spi_spi_control_port_write -> fpga_spi:write_n
	wire  [15:0] mm_interconnect_0_fpga_spi_spi_control_port_writedata;                       // mm_interconnect_0:fpga_spi_spi_control_port_writedata -> fpga_spi:data_from_cpu
	wire         mm_interconnect_0_dac_spi_spi_control_port_chipselect;                       // mm_interconnect_0:dac_spi_spi_control_port_chipselect -> dac_spi:spi_select
	wire  [15:0] mm_interconnect_0_dac_spi_spi_control_port_readdata;                         // dac_spi:data_to_cpu -> mm_interconnect_0:dac_spi_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_dac_spi_spi_control_port_address;                          // mm_interconnect_0:dac_spi_spi_control_port_address -> dac_spi:mem_addr
	wire         mm_interconnect_0_dac_spi_spi_control_port_read;                             // mm_interconnect_0:dac_spi_spi_control_port_read -> dac_spi:read_n
	wire         mm_interconnect_0_dac_spi_spi_control_port_write;                            // mm_interconnect_0:dac_spi_spi_control_port_write -> dac_spi:write_n
	wire  [15:0] mm_interconnect_0_dac_spi_spi_control_port_writedata;                        // mm_interconnect_0:dac_spi_spi_control_port_writedata -> dac_spi:data_from_cpu
	wire         mm_interconnect_0_flash_spi_spi_control_port_chipselect;                     // mm_interconnect_0:flash_spi_spi_control_port_chipselect -> flash_spi:spi_select
	wire  [15:0] mm_interconnect_0_flash_spi_spi_control_port_readdata;                       // flash_spi:data_to_cpu -> mm_interconnect_0:flash_spi_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_flash_spi_spi_control_port_address;                        // mm_interconnect_0:flash_spi_spi_control_port_address -> flash_spi:mem_addr
	wire         mm_interconnect_0_flash_spi_spi_control_port_read;                           // mm_interconnect_0:flash_spi_spi_control_port_read -> flash_spi:read_n
	wire         mm_interconnect_0_flash_spi_spi_control_port_write;                          // mm_interconnect_0:flash_spi_spi_control_port_write -> flash_spi:write_n
	wire  [15:0] mm_interconnect_0_flash_spi_spi_control_port_writedata;                      // mm_interconnect_0:flash_spi_spi_control_port_writedata -> flash_spi:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                                    // i2c_opencores_0:wb_inta_o -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                    // uart:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                    // fpga_spi:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                    // dac_spi:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                    // flash_spi:irq -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_cpu_irq_irq;                                                           // irq_mapper:sender_irq -> nios2_cpu:irq
	wire         rst_controller_reset_out_reset;                                              // rst_controller:reset_out -> [Av_FIFO_Int_0:rsi_nrst, dac_spi:reset_n, flash_spi:reset_n, fpga_spi:reset_n, i2c_opencores_0:wb_rst_i, irq_mapper:reset, leds:reset_n, lms_ctr_gpio:reset_n, mm_interconnect_0:nios2_cpu_reset_reset_bridge_in_reset_reset, nios2_cpu:reset_n, rst_translator:in_reset, switch:reset_n, sysid_qsys_0:reset_n, uart:reset_n]
	wire         rst_controller_reset_out_reset_req;                                          // rst_controller:reset_req -> [nios2_cpu:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                          // rst_controller_001:reset_out -> [dual_boot_0:nreset, mm_interconnect_0:dual_boot_0_nreset_reset_bridge_in_reset_reset, onchip_flash_0:reset_n, onchip_memory2_0:reset, rst_translator_001:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                                      // rst_controller_001:reset_req -> [onchip_memory2_0:reset_req, rst_translator_001:reset_req_in]

	avfifo #(
		.width (32)
	) av_fifo_int_0 (
		.clk            (clk_clk),                                                   //          clock.clk
		.address        (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect     (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_chipselect), //               .chipselect
		.write          (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_write),      //               .write
		.writedata      (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_writedata),  //               .writedata
		.read           (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_read),       //               .read
		.readdata       (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_readdata),   //               .readdata
		.rsi_nrst       (~rst_controller_reset_out_reset),                           //          reset.reset_n
		.coe_if_d       (exfifo_if_d_export),                                        //       cnd_if_d.export
		.coe_if_rd      (exfifo_if_rd_export),                                       //      cnd_if_rd.export
		.coe_of_wrfull  (exfifo_of_wrfull_export),                                   //  cnd_of_wrfull.export
		.coe_of_wr      (exfifo_of_wr_export),                                       //      cnd_of_wr.export
		.coe_of_d       (exfifo_of_d_export),                                        //       cnd_of_d.export
		.coe_if_rdempty (exfifo_if_rdempty_export),                                  // cnd_if_rdempty.export
		.coe_fifo_rst   (exfifo_rst_export)                                          //   cnd_fifo_rst.export
	);

	lms_ctr_dac_spi dac_spi (
		.clk           (clk_clk),                                               //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                       //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_dac_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_dac_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_dac_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_dac_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_dac_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_dac_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver3_irq),                              //              irq.irq
		.MISO          (dac_spi_ext_MISO),                                      //         external.export
		.MOSI          (dac_spi_ext_MOSI),                                      //                 .export
		.SCLK          (dac_spi_ext_SCLK),                                      //                 .export
		.SS_n          (dac_spi_ext_SS_n)                                       //                 .export
	);

	altera_dual_boot #(
		.INTENDED_DEVICE_FAMILY ("MAX 10"),
		.CONFIG_CYCLE           (15),
		.RESET_TIMER_CYCLE      (21)
	) dual_boot_0 (
		.clk                (clk_clk),                                        //    clk.clk
		.nreset             (~rst_controller_001_reset_out_reset),            // nreset.reset_n
		.avmm_rcv_address   (mm_interconnect_0_dual_boot_0_avalon_address),   // avalon.address
		.avmm_rcv_read      (mm_interconnect_0_dual_boot_0_avalon_read),      //       .read
		.avmm_rcv_writedata (mm_interconnect_0_dual_boot_0_avalon_writedata), //       .writedata
		.avmm_rcv_write     (mm_interconnect_0_dual_boot_0_avalon_write),     //       .write
		.avmm_rcv_readdata  (mm_interconnect_0_dual_boot_0_avalon_readdata)   //       .readdata
	);

	lms_ctr_flash_spi flash_spi (
		.clk           (clk_clk),                                                 //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                         //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_flash_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_flash_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_flash_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_flash_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_flash_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_flash_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver4_irq),                                //              irq.irq
		.MISO          (flash_spi_MISO),                                          //         external.export
		.MOSI          (flash_spi_MOSI),                                          //                 .export
		.SCLK          (flash_spi_SCLK),                                          //                 .export
		.SS_n          (flash_spi_SS_n)                                           //                 .export
	);

	lms_ctr_fpga_spi fpga_spi (
		.clk           (clk_clk),                                                //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                        //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_fpga_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_fpga_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_fpga_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_fpga_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_fpga_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_fpga_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver2_irq),                               //              irq.irq
		.MISO          (fpga_spi_ext_MISO),                                      //         external.export
		.MOSI          (fpga_spi_ext_MOSI),                                      //                 .export
		.SCLK          (fpga_spi_ext_SCLK),                                      //                 .export
		.SS_n          (fpga_spi_ext_SS_n)                                       //                 .export
	);

	i2c_opencores i2c_opencores_0 (
		.wb_clk_i   (clk_clk),                                                      //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                               //      clock_reset.reset
		.scl_pad_io (i2c_scl_export),                                               //       export_scl.export
		.sda_pad_io (i2c_sda_export),                                               //       export_sda.export
		.wb_adr_i   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver0_irq)                                      // interrupt_sender.irq
	);

	lms_ctr_leds leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_external_connection_export)       // external_connection.export
	);

	lms_ctr_lms_ctr_gpio lms_ctr_gpio (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_lms_ctr_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lms_ctr_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lms_ctr_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lms_ctr_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lms_ctr_gpio_s1_readdata),   //                    .readdata
		.out_port   (lms_ctr_gpio_external_connection_export)       // external_connection.export
	);

	lms_ctr_nios2_cpu nios2_cpu (
		.clk                                 (clk_clk),                                                 //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                         //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                      //                          .reset_req
		.d_address                           (nios2_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_cpu_data_master_read),                              //                          .read
		.d_readdata                          (nios2_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_cpu_data_master_write),                             //                          .write
		.d_writedata                         (nios2_cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),   //                          .writedata
		.E_ci_result                         (nios2_cpu_custom_instruction_master_result),              // custom_instruction_master.result
		.D_ci_a                              (nios2_cpu_custom_instruction_master_a),                   //                          .a
		.D_ci_b                              (nios2_cpu_custom_instruction_master_b),                   //                          .b
		.D_ci_c                              (nios2_cpu_custom_instruction_master_c),                   //                          .c
		.D_ci_n                              (nios2_cpu_custom_instruction_master_n),                   //                          .n
		.D_ci_readra                         (nios2_cpu_custom_instruction_master_readra),              //                          .readra
		.D_ci_readrb                         (nios2_cpu_custom_instruction_master_readrb),              //                          .readrb
		.D_ci_writerc                        (nios2_cpu_custom_instruction_master_writerc),             //                          .writerc
		.E_ci_dataa                          (nios2_cpu_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_datab                          (nios2_cpu_custom_instruction_master_datab),               //                          .datab
		.E_ci_multi_clock                    (),                                                        //                          .clk
		.E_ci_multi_reset                    (),                                                        //                          .reset
		.E_ci_multi_reset_req                (),                                                        //                          .reset_req
		.W_ci_estatus                        (nios2_cpu_custom_instruction_master_estatus),             //                          .estatus
		.W_ci_ipending                       (nios2_cpu_custom_instruction_master_ipending)             //                          .ipending
	);

	bitswap_qsys nios_custom_instr_bitswap_0 (
		.dataa  (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // s1.dataa
		.datab  (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //   .datab
		.result (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_result)  //   .result
	);

	altera_onchip_flash #(
		.INIT_FILENAME                       ("lms_ctr_onchip_flash_0.hex"),
		.INIT_FILENAME_SIM                   ("lms_ctr_onchip_flash_0.dat"),
		.DEVICE_FAMILY                       ("MAX 10"),
		.PART_NAME                           ("10M16SAU169C8G"),
		.DEVICE_ID                           ("16"),
		.SECTOR1_START_ADDR                  (0),
		.SECTOR1_END_ADDR                    (4095),
		.SECTOR2_START_ADDR                  (4096),
		.SECTOR2_END_ADDR                    (8191),
		.SECTOR3_START_ADDR                  (8192),
		.SECTOR3_END_ADDR                    (47103),
		.SECTOR4_START_ADDR                  (47104),
		.SECTOR4_END_ADDR                    (75775),
		.SECTOR5_START_ADDR                  (75776),
		.SECTOR5_END_ADDR                    (143359),
		.MIN_VALID_ADDR                      (0),
		.MAX_VALID_ADDR                      (143359),
		.MIN_UFM_VALID_ADDR                  (0),
		.MAX_UFM_VALID_ADDR                  (8191),
		.SECTOR1_MAP                         (1),
		.SECTOR2_MAP                         (2),
		.SECTOR3_MAP                         (3),
		.SECTOR4_MAP                         (4),
		.SECTOR5_MAP                         (5),
		.ADDR_RANGE1_END_ADDR                (143359),
		.ADDR_RANGE2_END_ADDR                (143359),
		.ADDR_RANGE1_OFFSET                  (1024),
		.ADDR_RANGE2_OFFSET                  (0),
		.ADDR_RANGE3_OFFSET                  (0),
		.AVMM_DATA_ADDR_WIDTH                (18),
		.AVMM_DATA_DATA_WIDTH                (32),
		.AVMM_DATA_BURSTCOUNT_WIDTH          (4),
		.SECTOR_READ_PROTECTION_MODE         (1),
		.FLASH_SEQ_READ_DATA_COUNT           (4),
		.FLASH_ADDR_ALIGNMENT_BITS           (2),
		.FLASH_READ_CYCLE_MAX_INDEX          (4),
		.FLASH_RESET_CYCLE_MAX_INDEX         (10),
		.FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  (48),
		.FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX (14000000),
		.FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX (12200),
		.PARALLEL_MODE                       (1),
		.READ_AND_WRITE_MODE                 (1),
		.WRAPPING_BURST_MODE                 (0),
		.IS_DUAL_BOOT                        ("True"),
		.IS_ERAM_SKIP                        ("True"),
		.IS_COMPRESSED_IMAGE                 ("True")
	) onchip_flash_0 (
		.clock                   (clk_clk),                                             //    clk.clk
		.reset_n                 (~rst_controller_001_reset_out_reset),                 // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_0_onchip_flash_0_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_0_onchip_flash_0_data_read),          //       .read
		.avmm_data_writedata     (mm_interconnect_0_onchip_flash_0_data_writedata),     //       .writedata
		.avmm_data_write         (mm_interconnect_0_onchip_flash_0_data_write),         //       .write
		.avmm_data_readdata      (mm_interconnect_0_onchip_flash_0_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_0_onchip_flash_0_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_0_onchip_flash_0_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_0_onchip_flash_0_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (mm_interconnect_0_onchip_flash_0_csr_address),        //    csr.address
		.avmm_csr_read           (mm_interconnect_0_onchip_flash_0_csr_read),           //       .read
		.avmm_csr_writedata      (mm_interconnect_0_onchip_flash_0_csr_writedata),      //       .writedata
		.avmm_csr_write          (mm_interconnect_0_onchip_flash_0_csr_write),          //       .write
		.avmm_csr_readdata       (mm_interconnect_0_onchip_flash_0_csr_readdata)        //       .readdata
	);

	lms_ctr_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	lms_ctr_switch switch (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_switch_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switch_s1_readdata), //                    .readdata
		.in_port  (switch_external_connection_export)     // external_connection.export
	);

	lms_ctr_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	lms_ctr_uart uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.rxd           (uart_external_connection_rxd),            // external_connection.export
		.txd           (uart_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver1_irq)                 //                 irq.irq
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) nios2_cpu_custom_instruction_master_translator (
		.ci_slave_dataa            (nios2_cpu_custom_instruction_master_dataa),                              //       ci_slave.dataa
		.ci_slave_datab            (nios2_cpu_custom_instruction_master_datab),                              //               .datab
		.ci_slave_result           (nios2_cpu_custom_instruction_master_result),                             //               .result
		.ci_slave_n                (nios2_cpu_custom_instruction_master_n),                                  //               .n
		.ci_slave_readra           (nios2_cpu_custom_instruction_master_readra),                             //               .readra
		.ci_slave_readrb           (nios2_cpu_custom_instruction_master_readrb),                             //               .readrb
		.ci_slave_writerc          (nios2_cpu_custom_instruction_master_writerc),                            //               .writerc
		.ci_slave_a                (nios2_cpu_custom_instruction_master_a),                                  //               .a
		.ci_slave_b                (nios2_cpu_custom_instruction_master_b),                                  //               .b
		.ci_slave_c                (nios2_cpu_custom_instruction_master_c),                                  //               .c
		.ci_slave_ipending         (nios2_cpu_custom_instruction_master_ipending),                           //               .ipending
		.ci_slave_estatus          (nios2_cpu_custom_instruction_master_estatus),                            //               .estatus
		.comb_ci_master_dataa      (nios2_cpu_custom_instruction_master_translator_comb_ci_master_dataa),    // comb_ci_master.dataa
		.comb_ci_master_datab      (nios2_cpu_custom_instruction_master_translator_comb_ci_master_datab),    //               .datab
		.comb_ci_master_result     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_result),   //               .result
		.comb_ci_master_n          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_n),        //               .n
		.comb_ci_master_readra     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_readra),   //               .readra
		.comb_ci_master_readrb     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_readrb),   //               .readrb
		.comb_ci_master_writerc    (nios2_cpu_custom_instruction_master_translator_comb_ci_master_writerc),  //               .writerc
		.comb_ci_master_a          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_a),        //               .a
		.comb_ci_master_b          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_b),        //               .b
		.comb_ci_master_c          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_c),        //               .c
		.comb_ci_master_ipending   (nios2_cpu_custom_instruction_master_translator_comb_ci_master_ipending), //               .ipending
		.comb_ci_master_estatus    (nios2_cpu_custom_instruction_master_translator_comb_ci_master_estatus),  //               .estatus
		.ci_slave_multi_clk        (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_reset      (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_clken      (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_reset_req  (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_start      (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_done       (),                                                                       //    (terminated)
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                   //    (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                   //    (terminated)
		.ci_slave_multi_result     (),                                                                       //    (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                            //    (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_a          (5'b00000),                                                               //    (terminated)
		.ci_slave_multi_b          (5'b00000),                                                               //    (terminated)
		.ci_slave_multi_c          (5'b00000),                                                               //    (terminated)
		.multi_ci_master_clk       (),                                                                       //    (terminated)
		.multi_ci_master_reset     (),                                                                       //    (terminated)
		.multi_ci_master_clken     (),                                                                       //    (terminated)
		.multi_ci_master_reset_req (),                                                                       //    (terminated)
		.multi_ci_master_start     (),                                                                       //    (terminated)
		.multi_ci_master_done      (1'b0),                                                                   //    (terminated)
		.multi_ci_master_dataa     (),                                                                       //    (terminated)
		.multi_ci_master_datab     (),                                                                       //    (terminated)
		.multi_ci_master_result    (32'b00000000000000000000000000000000),                                   //    (terminated)
		.multi_ci_master_n         (),                                                                       //    (terminated)
		.multi_ci_master_readra    (),                                                                       //    (terminated)
		.multi_ci_master_readrb    (),                                                                       //    (terminated)
		.multi_ci_master_writerc   (),                                                                       //    (terminated)
		.multi_ci_master_a         (),                                                                       //    (terminated)
		.multi_ci_master_b         (),                                                                       //    (terminated)
		.multi_ci_master_c         ()                                                                        //    (terminated)
	);

	lms_ctr_nios2_cpu_custom_instruction_master_comb_xconnect nios2_cpu_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (nios2_cpu_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (nios2_cpu_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (nios2_cpu_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (nios2_cpu_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (nios2_cpu_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (1)
	) nios2_cpu_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (),                                                                            // (terminated)
		.ci_master_readra    (),                                                                            // (terminated)
		.ci_master_readrb    (),                                                                            // (terminated)
		.ci_master_writerc   (),                                                                            // (terminated)
		.ci_master_a         (),                                                                            // (terminated)
		.ci_master_b         (),                                                                            // (terminated)
		.ci_master_c         (),                                                                            // (terminated)
		.ci_master_ipending  (),                                                                            // (terminated)
		.ci_master_estatus   (),                                                                            // (terminated)
		.ci_master_clk       (),                                                                            // (terminated)
		.ci_master_clken     (),                                                                            // (terminated)
		.ci_master_reset_req (),                                                                            // (terminated)
		.ci_master_reset     (),                                                                            // (terminated)
		.ci_master_start     (),                                                                            // (terminated)
		.ci_master_done      (1'b0),                                                                        // (terminated)
		.ci_slave_clk        (1'b0),                                                                        // (terminated)
		.ci_slave_clken      (1'b0),                                                                        // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                        // (terminated)
		.ci_slave_reset      (1'b0),                                                                        // (terminated)
		.ci_slave_start      (1'b0),                                                                        // (terminated)
		.ci_slave_done       ()                                                                             // (terminated)
	);

	lms_ctr_mm_interconnect_0 mm_interconnect_0 (
		.clk_main_clk_clk                               (clk_clk),                                                       //                             clk_main_clk.clk
		.dual_boot_0_nreset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                            // dual_boot_0_nreset_reset_bridge_in_reset.reset
		.nios2_cpu_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                                //    nios2_cpu_reset_reset_bridge_in_reset.reset
		.nios2_cpu_data_master_address                  (nios2_cpu_data_master_address),                                 //                    nios2_cpu_data_master.address
		.nios2_cpu_data_master_waitrequest              (nios2_cpu_data_master_waitrequest),                             //                                         .waitrequest
		.nios2_cpu_data_master_byteenable               (nios2_cpu_data_master_byteenable),                              //                                         .byteenable
		.nios2_cpu_data_master_read                     (nios2_cpu_data_master_read),                                    //                                         .read
		.nios2_cpu_data_master_readdata                 (nios2_cpu_data_master_readdata),                                //                                         .readdata
		.nios2_cpu_data_master_write                    (nios2_cpu_data_master_write),                                   //                                         .write
		.nios2_cpu_data_master_writedata                (nios2_cpu_data_master_writedata),                               //                                         .writedata
		.nios2_cpu_data_master_debugaccess              (nios2_cpu_data_master_debugaccess),                             //                                         .debugaccess
		.nios2_cpu_instruction_master_address           (nios2_cpu_instruction_master_address),                          //             nios2_cpu_instruction_master.address
		.nios2_cpu_instruction_master_waitrequest       (nios2_cpu_instruction_master_waitrequest),                      //                                         .waitrequest
		.nios2_cpu_instruction_master_read              (nios2_cpu_instruction_master_read),                             //                                         .read
		.nios2_cpu_instruction_master_readdata          (nios2_cpu_instruction_master_readdata),                         //                                         .readdata
		.Av_FIFO_Int_0_avalon_slave_0_address           (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_address),        //             Av_FIFO_Int_0_avalon_slave_0.address
		.Av_FIFO_Int_0_avalon_slave_0_write             (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_write),          //                                         .write
		.Av_FIFO_Int_0_avalon_slave_0_read              (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_read),           //                                         .read
		.Av_FIFO_Int_0_avalon_slave_0_readdata          (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_readdata),       //                                         .readdata
		.Av_FIFO_Int_0_avalon_slave_0_writedata         (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_writedata),      //                                         .writedata
		.Av_FIFO_Int_0_avalon_slave_0_chipselect        (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_chipselect),     //                                         .chipselect
		.dac_spi_spi_control_port_address               (mm_interconnect_0_dac_spi_spi_control_port_address),            //                 dac_spi_spi_control_port.address
		.dac_spi_spi_control_port_write                 (mm_interconnect_0_dac_spi_spi_control_port_write),              //                                         .write
		.dac_spi_spi_control_port_read                  (mm_interconnect_0_dac_spi_spi_control_port_read),               //                                         .read
		.dac_spi_spi_control_port_readdata              (mm_interconnect_0_dac_spi_spi_control_port_readdata),           //                                         .readdata
		.dac_spi_spi_control_port_writedata             (mm_interconnect_0_dac_spi_spi_control_port_writedata),          //                                         .writedata
		.dac_spi_spi_control_port_chipselect            (mm_interconnect_0_dac_spi_spi_control_port_chipselect),         //                                         .chipselect
		.dual_boot_0_avalon_address                     (mm_interconnect_0_dual_boot_0_avalon_address),                  //                       dual_boot_0_avalon.address
		.dual_boot_0_avalon_write                       (mm_interconnect_0_dual_boot_0_avalon_write),                    //                                         .write
		.dual_boot_0_avalon_read                        (mm_interconnect_0_dual_boot_0_avalon_read),                     //                                         .read
		.dual_boot_0_avalon_readdata                    (mm_interconnect_0_dual_boot_0_avalon_readdata),                 //                                         .readdata
		.dual_boot_0_avalon_writedata                   (mm_interconnect_0_dual_boot_0_avalon_writedata),                //                                         .writedata
		.flash_spi_spi_control_port_address             (mm_interconnect_0_flash_spi_spi_control_port_address),          //               flash_spi_spi_control_port.address
		.flash_spi_spi_control_port_write               (mm_interconnect_0_flash_spi_spi_control_port_write),            //                                         .write
		.flash_spi_spi_control_port_read                (mm_interconnect_0_flash_spi_spi_control_port_read),             //                                         .read
		.flash_spi_spi_control_port_readdata            (mm_interconnect_0_flash_spi_spi_control_port_readdata),         //                                         .readdata
		.flash_spi_spi_control_port_writedata           (mm_interconnect_0_flash_spi_spi_control_port_writedata),        //                                         .writedata
		.flash_spi_spi_control_port_chipselect          (mm_interconnect_0_flash_spi_spi_control_port_chipselect),       //                                         .chipselect
		.fpga_spi_spi_control_port_address              (mm_interconnect_0_fpga_spi_spi_control_port_address),           //                fpga_spi_spi_control_port.address
		.fpga_spi_spi_control_port_write                (mm_interconnect_0_fpga_spi_spi_control_port_write),             //                                         .write
		.fpga_spi_spi_control_port_read                 (mm_interconnect_0_fpga_spi_spi_control_port_read),              //                                         .read
		.fpga_spi_spi_control_port_readdata             (mm_interconnect_0_fpga_spi_spi_control_port_readdata),          //                                         .readdata
		.fpga_spi_spi_control_port_writedata            (mm_interconnect_0_fpga_spi_spi_control_port_writedata),         //                                         .writedata
		.fpga_spi_spi_control_port_chipselect           (mm_interconnect_0_fpga_spi_spi_control_port_chipselect),        //                                         .chipselect
		.i2c_opencores_0_avalon_slave_0_address         (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address),      //           i2c_opencores_0_avalon_slave_0.address
		.i2c_opencores_0_avalon_slave_0_write           (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write),        //                                         .write
		.i2c_opencores_0_avalon_slave_0_readdata        (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata),     //                                         .readdata
		.i2c_opencores_0_avalon_slave_0_writedata       (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata),    //                                         .writedata
		.i2c_opencores_0_avalon_slave_0_waitrequest     (~mm_interconnect_0_i2c_opencores_0_avalon_slave_0_waitrequest), //                                         .waitrequest
		.i2c_opencores_0_avalon_slave_0_chipselect      (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect),   //                                         .chipselect
		.leds_s1_address                                (mm_interconnect_0_leds_s1_address),                             //                                  leds_s1.address
		.leds_s1_write                                  (mm_interconnect_0_leds_s1_write),                               //                                         .write
		.leds_s1_readdata                               (mm_interconnect_0_leds_s1_readdata),                            //                                         .readdata
		.leds_s1_writedata                              (mm_interconnect_0_leds_s1_writedata),                           //                                         .writedata
		.leds_s1_chipselect                             (mm_interconnect_0_leds_s1_chipselect),                          //                                         .chipselect
		.lms_ctr_gpio_s1_address                        (mm_interconnect_0_lms_ctr_gpio_s1_address),                     //                          lms_ctr_gpio_s1.address
		.lms_ctr_gpio_s1_write                          (mm_interconnect_0_lms_ctr_gpio_s1_write),                       //                                         .write
		.lms_ctr_gpio_s1_readdata                       (mm_interconnect_0_lms_ctr_gpio_s1_readdata),                    //                                         .readdata
		.lms_ctr_gpio_s1_writedata                      (mm_interconnect_0_lms_ctr_gpio_s1_writedata),                   //                                         .writedata
		.lms_ctr_gpio_s1_chipselect                     (mm_interconnect_0_lms_ctr_gpio_s1_chipselect),                  //                                         .chipselect
		.nios2_cpu_debug_mem_slave_address              (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),           //                nios2_cpu_debug_mem_slave.address
		.nios2_cpu_debug_mem_slave_write                (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),             //                                         .write
		.nios2_cpu_debug_mem_slave_read                 (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),              //                                         .read
		.nios2_cpu_debug_mem_slave_readdata             (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),          //                                         .readdata
		.nios2_cpu_debug_mem_slave_writedata            (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),         //                                         .writedata
		.nios2_cpu_debug_mem_slave_byteenable           (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),        //                                         .byteenable
		.nios2_cpu_debug_mem_slave_waitrequest          (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest),       //                                         .waitrequest
		.nios2_cpu_debug_mem_slave_debugaccess          (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess),       //                                         .debugaccess
		.onchip_flash_0_csr_address                     (mm_interconnect_0_onchip_flash_0_csr_address),                  //                       onchip_flash_0_csr.address
		.onchip_flash_0_csr_write                       (mm_interconnect_0_onchip_flash_0_csr_write),                    //                                         .write
		.onchip_flash_0_csr_read                        (mm_interconnect_0_onchip_flash_0_csr_read),                     //                                         .read
		.onchip_flash_0_csr_readdata                    (mm_interconnect_0_onchip_flash_0_csr_readdata),                 //                                         .readdata
		.onchip_flash_0_csr_writedata                   (mm_interconnect_0_onchip_flash_0_csr_writedata),                //                                         .writedata
		.onchip_flash_0_data_address                    (mm_interconnect_0_onchip_flash_0_data_address),                 //                      onchip_flash_0_data.address
		.onchip_flash_0_data_write                      (mm_interconnect_0_onchip_flash_0_data_write),                   //                                         .write
		.onchip_flash_0_data_read                       (mm_interconnect_0_onchip_flash_0_data_read),                    //                                         .read
		.onchip_flash_0_data_readdata                   (mm_interconnect_0_onchip_flash_0_data_readdata),                //                                         .readdata
		.onchip_flash_0_data_writedata                  (mm_interconnect_0_onchip_flash_0_data_writedata),               //                                         .writedata
		.onchip_flash_0_data_burstcount                 (mm_interconnect_0_onchip_flash_0_data_burstcount),              //                                         .burstcount
		.onchip_flash_0_data_readdatavalid              (mm_interconnect_0_onchip_flash_0_data_readdatavalid),           //                                         .readdatavalid
		.onchip_flash_0_data_waitrequest                (mm_interconnect_0_onchip_flash_0_data_waitrequest),             //                                         .waitrequest
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),                 //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                   //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),                //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),               //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),              //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),              //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                   //                                         .clken
		.switch_s1_address                              (mm_interconnect_0_switch_s1_address),                           //                                switch_s1.address
		.switch_s1_readdata                             (mm_interconnect_0_switch_s1_readdata),                          //                                         .readdata
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),          //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),         //                                         .readdata
		.uart_s1_address                                (mm_interconnect_0_uart_s1_address),                             //                                  uart_s1.address
		.uart_s1_write                                  (mm_interconnect_0_uart_s1_write),                               //                                         .write
		.uart_s1_read                                   (mm_interconnect_0_uart_s1_read),                                //                                         .read
		.uart_s1_readdata                               (mm_interconnect_0_uart_s1_readdata),                            //                                         .readdata
		.uart_s1_writedata                              (mm_interconnect_0_uart_s1_writedata),                           //                                         .writedata
		.uart_s1_begintransfer                          (mm_interconnect_0_uart_s1_begintransfer),                       //                                         .begintransfer
		.uart_s1_chipselect                             (mm_interconnect_0_uart_s1_chipselect)                           //                                         .chipselect
	);

	lms_ctr_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (nios2_cpu_irq_irq)               //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_cpu_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_cpu_debug_reset_request_reset),    // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
